library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CU is port(
    clk, rst, interrupt, restart: in std_logic;
    instruction: in std_logic_vector(15 downto 0);
    jump_enable, jump_zero_enable, flag_feedback, mem_read_enable, pc_immediate,pc_write, restart_out, interrupt_out, push_flags, mem_write, is_in_port, is_immediate, stall_Fenable, stall_Eenable, stall_Menable, flag_enable, alu_mem, WB1_enable, WB2_enable, SP_enable, SP_op, SP_select,FB_enable, FB_op, outport_enable: out std_logic;
    WB1_addr, WB2_addr: out std_logic_vector(2 downto 0);
    alu_op: out std_logic_vector(3 downto 0)
);
end entity;

architecture Behavioral of CU is
TYPE state_type is(standards, NOP, interrupt_state, restart_state, return_state, RTI_state);
signal status: state_type := standards;
begin
    process(instruction, clk, rst, interrupt, restart)
    variable loaded_addr: std_logic_vector(2 downto 0);
    variable interrupt_cycles: integer := 0;
    variable restart_cycles: integer := 0;
    variable return_cycles: integer := 0;
    variable RTI_cycles: integer := 0;
    variable pop_hazard: std_logic := '0';
    variable true_stall: std_logic := '0';
    begin 
        if rst = '1' then
            status <= standards;
            WB1_enable <= '0';
            WB2_enable <= '0';
            is_in_port <= '0';
            is_immediate <= '0';
            stall_Fenable <= '0';
            stall_Eenable <= '0';
            flag_enable <= '0';
            mem_write <= '0';
            SP_enable <= '0';
            interrupt_out <= '0';
            outport_enable <= '0';
            FB_enable <= '0';
            alu_mem <= '0';
            alu_op <= "0000";
            pc_immediate <= '0';
            restart_out <= '0';
            push_flags <= '0';
            jump_enable <= '0';
            jump_zero_enable <= '0';
            mem_read_enable <= '0';
            flag_feedback <= '0';
        elsif interrupt = '1' then
            status <= interrupt_state;
            interrupt_cycles := 1;
            stall_Fenable <= '1';
            stall_Eenable <= '0';
            Wb1_enable <= '0';
            WB2_enable <= '0';
            is_in_port <= '0';
            is_immediate <= '1';
            flag_enable <= '0';
            mem_write <= '1';
            SP_enable <= '1';
            SP_op <= '1';
            SP_select <= '0';
            outport_enable <= '0';
            FB_enable <= '0';
            interrupt_out <= '1';
            alu_mem <= '1';
            alu_op <= "1101";
            pc_immediate <= '1';
            restart_out <= '0';
            push_flags <= '0';
            pc_write <= '1';
            jump_enable <= '0';
            jump_zero_enable <= '0';
            mem_read_enable <= '1';
            flag_feedback <= '0';
        elsif restart = '1' then
            status <= restart_state;
            restart_cycles := 1;
            WB1_enable <= '0';
            WB2_enable <= '0';
            is_in_port <= '0';
            is_immediate <= '0';
            stall_Fenable <= '1';
            flag_enable <= '0';
            interrupt_out <= '0';
            mem_write <= '0';
            SP_enable <= '0';
            pc_write <= '0';
            outport_enable <= '0';
            FB_enable <= '0';
            alu_mem <= '0';
            alu_op <= "1101";
            pc_immediate <= '1';
            push_flags <= '0';
            mem_read_enable <= '1';
            restart_out <= '1';
            jump_enable <= '0';
            jump_zero_enable <= '0';
            flag_feedback <= '0';
        else
            case status is
                when standards =>
                    restart_out <= '0';
                    interrupt_out <= '0';
                    flag_feedback <= '0';
                    stall_Menable <= '0';
                    if true_stall = '1' then
                        stall_Fenable <= '0';
                        stall_Eenable <= '0';
                        true_stall := '0';
                    end if;
                    if pop_hazard = '1' then
                        if instruction(15 downto 14) = "10" then
                            if loaded_addr = instruction(9 downto 7) or loaded_addr = instruction(6 downto 4) then
                                stall_Fenable <= '1';
                                true_stall := '1';
                            else
                            end if;
                        elsif instruction(15 downto 12) = "0100" then
                            if loaded_addr = instruction(9 downto 7) then
                                stall_Fenable <= '1';
                                true_stall := '1';
                            end if;
                        elsif not (instruction(15 downto 10) = "000111" or instruction(15 downto 10) = "000101") then
                            if loaded_addr = instruction(9 downto 7) then
                                stall_Fenable <= '1';
                                true_stall := '1';
                            end if;
                        else
                            null;
                        end if;
                        pop_hazard := '0';
                        loaded_addr := "000";
                    end if;
                    if true_stall = '0' then
                    case instruction(15 downto 10) is
                        when "100000" | "100001" | "100010" | "100011" | "100100"=>
                            WB1_enable <= '1';
                            WB1_addr <= instruction(3 downto 1);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '1';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            push_flags <= '0';
                            pc_write <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '0';
                        when "000001" | "000010" | "000011" | "000100" =>
                            WB1_enable <= '1';
                            WB1_addr <= instruction(9 downto 7);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '1';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            push_flags <= '0';
                            pc_immediate <= '0';
                            pc_write <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '0';
                        when "010000" | "010001" =>
                            wb1_enable <= '1';
                            wb1_addr <= instruction(3 downto 1);
                            wb2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '1';
                            flag_enable <= '1';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            push_flags <= '0';
                            alu_mem <= '0';
                            FB_enable <= '0';
                            pc_write <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            status <= NOP;
                            mem_read_enable <= '0';
                        when "010010" =>
                            status <= NOP;
                            WB1_enable <= '1';
                            WB1_addr <= instruction(3 downto 1);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '1';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '1';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            push_flags <= '0';
                            pc_write <= '0';
                            mem_read_enable <= '1';
                        when "010011" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '1';
                            flag_enable <= '0';
                            mem_write <= '1';
                            SP_enable <= '0';
                            SP_select <= '1';
                            outport_enable <= '0';
                            push_flags <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            pc_write <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            status <= NOP;
                            mem_read_enable <= '0';
                        when "100101" =>
                            WB1_enable <= '1';
                            WB1_addr <= instruction(3 downto 1);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            push_flags <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            pc_write <= '0';
                            alu_mem <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '1';
                        when "101001" =>
                            WB1_enable <= '1';
                            WB1_addr <= instruction(6 downto 4);
                            WB2_enable <= '1';
                            WB2_addr <= instruction(9 downto 7);
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            pc_write <= '0';
                            alu_mem <= '0';
                            push_flags <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '1';
                        when "101010" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '1';
                            push_flags <= '0';
                            mem_write <= '0';
                            alu_mem <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            pc_write <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '1';
                        when "000101" =>
                            WB1_enable <= '1';
                            WB1_addr <= instruction(9 downto 7);
                            WB2_enable <= '0';
                            is_in_port <= '1';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            pc_write <= '0';
                            SP_enable <= '0';
                            alu_mem <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            push_flags <= '0';
                            mem_read_enable <= '0';
                            jump_zero_enable <= '0';
                        when "000110" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            alu_mem <= '0';
                            outport_enable <= '1';
                            push_flags <= '0';
                            FB_enable <= '0';
                            pc_write <= '0';
                            mem_read_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "000111" =>
                            WB1_enable <= '1';
                            stall_Fenable <= '0';
                            loaded_addr := instruction(9 downto 7);
                            pop_hazard := '1';
                            stall_Eenable <= '0';
                            WB1_addr <= instruction(9 downto 7);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '1';
                            push_flags <= '0';
                            SP_enable <= '1';
                            SP_op <= '0';
                            SP_select <= '0';
                            mem_read_enable <= '1';
                            pc_write <= '0';
                            alu_mem <= '1';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "001000" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_read_enable <= '0';
                            push_flags <= '0';
                            mem_write <= '1';
                            SP_enable <= '1';
                            SP_op <= '1';
                            SP_select <= '0';
                            alu_mem <= '0';
                            pc_write <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "001001" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            push_flags <= '0';
                            SP_enable <= '0';
                            SP_select <= '0';
                            pc_write <= '0';
                            alu_mem <= '0';
                            outport_enable <= '0';
                            FB_enable <= '1';
                            FB_op <= '1';
                            mem_read_enable <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "001010" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            push_flags <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            SP_select <= '0';
                            alu_mem <= '0';
                            outport_enable <= '0';
                            FB_enable <= '1';
                            pc_write <= '0';
                            FB_op <= '0';
                            pc_immediate <= '0';
                            mem_read_enable <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "000000" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            alu_mem <= '0';
                            push_flags <= '0';
                            SP_enable <= '0';
                            pc_write <= '0';
                            outport_enable <= '0';
                            FB_enable <= '1';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                        when "010100" =>
                            status <= NOP;
                            WB1_enable <= '1';
                            WB1_addr <= instruction(3 downto 1);
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '1';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            pc_write <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            push_flags <= '0';
                            mem_read_enable <= '0';
                        when "110001" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            pc_write <= '0';
                            push_flags <= '0';
                            jump_enable <= '1';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '0';
                        when "110000" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '0';
                            outport_enable <= '0';
                            push_flags <= '0';
                            pc_write <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '1';
                            mem_read_enable <= '0';
                        when "110010" =>
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '1';
                            flag_enable <= '0';
                            mem_write <= '1';
                            SP_enable <= '1';
                            Sp_op <= '1';
                            SP_select <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '1';
                            push_flags <= '0';
                            pc_write <= '0';
                            jump_enable <= '1';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '0';
                        when "110011" =>
                            status <= return_state;
                            stall_Fenable <= '1';
                            stall_Eenable <= '0';
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '1';
                            SP_op <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            push_flags <= '0';
                            pc_write <= '1';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '1';
                            return_cycles := 1;
                        when "110100" =>
                            status <= RTI_state;
                            stall_Fenable <= '1';
                            stall_Eenable <= '0';
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            SP_enable <= '1';
                            SP_op <= '0';
                            sp_select <= '0';
                            outport_enable <= '0';
                            flag_feedback <= '1';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            pc_immediate <= '0';
                            push_flags <= '0';
                            pc_write <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '1';
                            RTI_cycles := 1;
                        when others =>
                            null;
                        end case;
                        case instruction(15 downto 10) is
                            when "100000" | "010000" | "010011" | "010010"=> alu_op <= "1000";
                            when "100001" | "010001" => alu_op <= "1001";
                            when "100010" => alu_op <= "0010";
                            when "100011" => alu_op <= "0011";
                            when "100100" => alu_op <= "0100";
                            when "010100" | "110010" => alu_op <= "0001";
                            when "101010" => alu_op <= "0110";
                            when "000001" => alu_op <= "0101";
                            when "000010" => alu_op <= "1100";
                            when "000011" => alu_op <= "1010";
                            when "000100" => alu_op <= "1011";
                            when "000111" | "110100" => alu_op <= "1111";
                            when others => alu_op <= "0000";
                        end case;
                    else
                        wb1_enable <= '0';
                        wb2_enable <= '0';
                        is_in_port <= '0';
                        is_immediate <= '0';
                        flag_enable <= '0';
                        mem_write <= '0';
                        SP_enable <= '0';
                        outport_enable <= '0';
                        FB_enable <= '0';
                        alu_mem <= '0';
                        pc_immediate <= '0';
                        push_flags <= '0';
                        pc_write <= '0';
                        jump_enable <= '0';
                        jump_zero_enable <= '0';
                        mem_read_enable <= '0';
                        alu_op <= "0000";
                    end if;
                when NOP => 
                    stall_Fenable <= '0';
                    stall_Eenable <= '0';
                    WB1_enable <= '0';
                    WB2_enable <= '0';
                    is_in_port <= '0';
                    is_immediate <= '0';
                    flag_enable <= '0';
                    mem_write <= '0';
                    push_flags <= '0';
                    alu_mem <= '0';
                    SP_enable <= '0';
                    outport_enable <= '0';
                    FB_enable <= '0';
                    pc_immediate <= '0';
                    interrupt_out <= '0';
                    pc_write <= '0';
                    mem_read_enable <= '0';
                    alu_op <= "0001";
                    status <= standards;
                when RTI_state =>
                    if RTI_cycles < 4 then
                        if RTI_cycles = 1 then
                            flag_feedback <= '0';
                            pc_write <= '1';
                        else
                            interrupt_out <= '0';
                            stall_Eenable <= '0';
                            flag_feedback <= '0';
                            SP_enable <= '0';
                            SP_op <= '0';
                            pc_write <= '0';
                            push_flags <= '0';
                            pc_immediate <= '0';
                            WB1_enable <= '0';
                            WB2_enable <= '0';
                            is_in_port <= '0';
                            is_immediate <= '0';
                            flag_enable <= '0';
                            mem_write <= '0';
                            outport_enable <= '0';
                            FB_enable <= '0';
                            alu_mem <= '0';
                            jump_enable <= '0';
                            jump_zero_enable <= '0';
                            mem_read_enable <= '0';
                        end if;
                        RTI_cycles := RTI_cycles + 1;
                        stall_Fenable <= '1';
                    else
                        RTI_cycles := 0;
                        mem_read_enable <= '0';
                        stall_Fenable <= '0';
                        stall_Eenable <= '0';
                        pc_write <= '0';
                        SP_enable <= '0';
                        status <= standards;
                    end if;
                when return_state =>
                    if return_cycles < 4 then
                        WB1_enable <= '0';
                        WB2_enable <= '0';
                        is_in_port <= '0';
                        is_immediate <= '0';
                        flag_enable <= '0';
                        mem_write <= '0';
                        SP_enable <= '0';
                        outport_enable <= '0';
                        FB_enable <= '0';
                        alu_mem <= '0';
                        pc_immediate <= '0';
                        push_flags <= '0';
                        pc_write <= '0';
                        jump_enable <= '0';
                        jump_zero_enable <= '0';
                        mem_read_enable <= '0';
                        return_cycles := return_cycles + 1;
                        stall_Fenable <= '1';
                    else
                        return_cycles := 0;
                        stall_Fenable <= '0';
                        stall_Eenable <= '0';
                        status <= standards;
                    end if;
                when interrupt_state =>
                    if interrupt_cycles < 3 then
                        if interrupt_cycles = 1 then
                            push_flags <= '1';
                            interrupt_out <= '0';
                            stall_Fenable <= '1';
                            stall_Eenable <= '0';
                            pc_write <= '0';
                        else
                            push_flags <= '0';
                            SP_enable <= '0';
                            pc_immediate <= '0';
                            stall_Fenable <= '1';
                            stall_Eenable <= '1';
                        end if;
                        interrupt_cycles := interrupt_cycles + 1;
                    else
                        interrupt_cycles := 0;
                        stall_Fenable <= '0';
                        stall_eenable <= '0';
                        status <= standards;
                    end if;
                when restart_state =>
                    if restart_cycles < 3 then
                        restart_cycles := restart_cycles + 1;
                        stall_Fenable <= '1';
                        stall_Eenable <= '1';
                    else
                        restart_cycles := 0;
                        stall_Fenable <= '0';
                        stall_Eenable <= '0';
                        status <= standards;
                    end if;
                    restart_out <= '0';
            end case;
        end if;
    end process;
end architecture;